module game_process(
    matrix_out,
    x_pos,
    y_pos,
    player_top,
    player_down,
    count,
    clk
);

parameter SIZE = 2;
parameter WIDTH = 8;
parameter BIT_OF_WIDTH = 3;

output[15:0] matrix_out;
reg[15:0] matrix_out;

input[2:0] player_top, player_down;

input[BIT_OF_WIDTH-1:0] x_pos, y_pos;

input clk;
input[2:0] count;

integer i;

always @ (posedge clk)
begin
	matrix_out = 0;
    // top player
	if(count == 0)begin
        case(player_top)
            0 : matrix_out = 8'b00000011; 
            1 : matrix_out = 8'b00000110; 
            2 : matrix_out = 8'b00001100; 
            3 : matrix_out = 8'b00011000; 
            4 : matrix_out = 8'b00110000; 
            5 : matrix_out = 8'b01100000; 
            6 : matrix_out = 8'b11000000; 
            7 : matrix_out = 0;
        endcase
	end
    // down player
	if(count == 7)begin
        case (player_down)
            0 : matrix_out = 8'b00000011; 
            1 : matrix_out = 8'b00000110; 
            2 : matrix_out = 8'b00001100; 
            3 : matrix_out = 8'b00011000; 
            4 : matrix_out = 8'b00110000; 
            5 : matrix_out = 8'b01100000; 
            6 : matrix_out = 8'b11000000; 
			7 : matrix_out = 0;
        endcase
	end
	// ball
    if(count == y_pos) begin
        for(i = 0; i < WIDTH; i = i + 1) begin
            matrix_out[i] = (x_pos == i) ? 1 : matrix_out[i];
        end
    end
end

endmodule // game_process
