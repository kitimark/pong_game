module testtt(
    in,
    out
);

input[2:0] in;
output[2:0] out;

assign out = in;

endmodule // testtt